--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   16:23:59 04/01/2024
-- Design Name:   
-- Module Name:   /home/student/Desktop/13000122098/one_to_eight_demux/one_to_eight_demux_test.vhd
-- Project Name:  one_to_eight_demux
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: one_to_eight_demux_rtl
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY one_to_eight_demux_test IS
END one_to_eight_demux_test;
 
ARCHITECTURE behavior OF one_to_eight_demux_test IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT one_to_eight_demux_rtl
    PORT(
         d : IN  std_logic;
         s : IN  std_logic_vector(2 downto 0);
         o : OUT  std_logic_vector(7 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal d : std_logic := '0';
   signal s : std_logic_vector(2 downto 0) := (others => '0');

 	--Outputs
   signal o : std_logic_vector(7 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
 
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: one_to_eight_demux_rtl PORT MAP (
          d => d,
          s => s,
          o => o
        );

   -- Clock process definitions

 

   -- Stimulus process
   stim_proc: process
   begin		
     d<='1';
	  s<="000";
	  wait for 1 ps;
	  d<='1';
	  s<="001";
	  wait for 1 ps;
	  d<='1';
	  s<="010";
	  wait for 1 ps;
	  d<='1';
	  s<="011";
	  wait for 1 ps;
	  d<='1';
	  s<="100";
	  wait for 1 ps;
	  d<='1';
	  s<="101";
	  wait for 1 ps;
	  d<='1';
	  s<="110";
	  wait for 1 ps;
	  d<='1';
	  s<="111";
	  wait for 1 ps;
   end process;

END;
